Name 19----/19d----,resistive transient analysis

**parameter 
.temp 27 

**input 
vin 1 0 sin(0 1 1k)


**circuit 
r1 1 2 1k
r2 2 0 1k 
r3 2 3 1k 
r4 3 0 1k

**command 
.tran 0.1m 1m 

.end 
